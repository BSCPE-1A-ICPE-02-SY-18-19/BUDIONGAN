CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
140 0 18 100 10
214 107 1172 613
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
382 203 495 300
9437202 0
0
6 Title:
5 Name:
0
0
0
10
7 Pulser~
4 202 208 0 10 12
0 17 18 19 15 0 0 5 5 5
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
7168 0 0
2
43530.4 0
0
2 +V
167 299 67 0 1 3
0 3
0
0 0 54256 0
3 10V
-9 -22 12 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3171 0 0
2
43530.4 0
0
6 74LS48
188 814 131 0 14 29
0 14 2 6 4 20 21 7 8 9
10 11 12 13 22
0
0 0 4848 0
7 74LS248
-24 -60 25 -52
2 U5
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 0 0 0 0
1 U
4139 0 0
2
43530.3 0
0
9 CC 7-Seg~
183 972 133 0 18 19
10 13 12 11 10 9 8 7 23 24
0 0 0 1 1 1 1 2 2
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
6435 0 0
2
5.89883e-315 0
0
6 74112~
219 530 165 0 7 32
0 3 5 15 5 3 25 2
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U4A
-30 2 -9 10
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 4 0
1 U
5283 0 0
2
5.89883e-315 0
0
9 2-In AND~
219 576 60 0 3 22
0 5 2 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -5 9 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
6874 0 0
2
5.89883e-315 0
0
9 2-In AND~
219 485 51 0 3 22
0 4 6 5
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-14 -5 7 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5305 0 0
2
5.89883e-315 0
0
6 74112~
219 645 165 0 7 32
0 3 16 15 16 3 26 14
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
-26 1 -5 9
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
34 0 0
2
5.89883e-315 0
0
6 74112~
219 415 164 0 7 32
0 3 4 15 4 3 27 6
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1B
-27 1 -6 9
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
969 0 0
2
5.89883e-315 0
0
6 74112~
219 299 164 0 7 32
0 3 28 15 29 3 30 4
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1A
-29 1 -8 9
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
8402 0 0
2
5.89883e-315 0
0
35
0 2 2 0 0 4224 0 0 3 33 0 4
554 92
742 92
742 104
782 104
0 0 3 0 0 4096 0 0 0 15 13 2
576 102
576 177
0 0 3 0 0 0 0 0 0 14 12 2
461 102
461 176
0 0 3 0 0 0 0 0 0 16 11 2
357 101
357 176
0 1 4 0 0 8192 0 0 7 6 0 3
370 128
370 42
461 42
4 0 4 0 0 0 0 9 0 0 35 3
391 146
370 146
370 128
1 1 3 0 0 0 0 10 2 0 0 2
299 101
299 76
0 0 5 0 0 4224 0 0 0 31 32 3
492 129
492 69
518 69
0 4 4 0 0 8320 0 0 3 35 0 5
334 128
334 226
766 226
766 122
782 122
0 3 6 0 0 12416 0 0 3 34 0 6
439 119
450 119
450 217
758 217
758 113
782 113
5 5 3 0 0 4224 0 9 10 0 0 2
415 176
299 176
5 5 3 0 0 0 0 5 9 0 0 3
530 177
530 176
415 176
5 5 3 0 0 0 0 8 5 0 0 2
645 177
530 177
1 1 3 0 0 0 0 9 5 0 0 3
415 101
415 102
530 102
1 1 3 0 0 0 0 5 8 0 0 2
530 102
645 102
1 1 3 0 0 128 0 10 9 0 0 2
299 101
415 101
7 7 7 0 0 8320 0 3 4 0 0 5
846 95
912 95
912 207
987 207
987 169
8 6 8 0 0 8320 0 3 4 0 0 5
846 104
917 104
917 202
981 202
981 169
9 5 9 0 0 8320 0 3 4 0 0 5
846 113
922 113
922 197
975 197
975 169
10 4 10 0 0 4224 0 3 4 0 0 5
846 122
927 122
927 192
969 192
969 169
11 3 11 0 0 4224 0 3 4 0 0 5
846 131
932 131
932 187
963 187
963 169
12 2 12 0 0 4224 0 3 4 0 0 5
846 140
937 140
937 182
957 182
957 169
13 1 13 0 0 4224 0 3 4 0 0 5
846 149
942 149
942 177
951 177
951 169
7 1 14 0 0 4224 0 8 3 0 0 4
669 129
749 129
749 95
782 95
3 0 15 0 0 8192 0 5 0 0 28 3
500 138
473 138
473 208
3 0 15 0 0 8192 0 9 0 0 28 3
385 137
381 137
381 208
3 0 15 0 0 0 0 10 0 0 28 3
269 137
254 137
254 208
4 3 15 0 0 4224 0 1 8 0 0 4
232 208
608 208
608 138
615 138
0 2 16 0 0 4096 0 0 8 30 0 2
598 129
621 129
3 4 16 0 0 4224 0 6 8 0 0 5
597 60
597 104
598 104
598 147
621 147
2 4 5 0 0 0 0 5 5 0 0 6
506 129
492 129
492 131
491 131
491 147
506 147
3 1 5 0 0 128 0 7 6 0 0 6
506 51
518 51
518 69
518 69
518 51
552 51
7 2 2 0 0 128 0 5 6 0 0 3
554 129
554 69
552 69
7 2 6 0 0 128 0 9 7 0 0 3
439 128
439 60
461 60
7 2 4 0 0 128 0 10 9 0 0 2
323 128
391 128
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
